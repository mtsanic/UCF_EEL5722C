`timescale 1ns / 1ps


module pause_rom(
        input wire clk,
        input wire pause,
		input wire [9:0] x,
		input wire [9:0] y,
        output pause_on,
		output [11:0] pause_rgb
);

(* rom_style = "block" *)

    localparam  X_START = 263,
                X_END   = 361,
                Y_START = 206,
                Y_END   = 224;

    reg [3:0] rows;
    reg [6:0] cols;
    reg  b_rgb;

    always @(posedge clk)
		begin
		rows <= y - Y_START - 1;
		cols <= x - X_START - 1;
		end
    
    always @(*) begin
            case ({cols,rows})

                // P character

                11'b000_0100_0011 : b_rgb<=1'b1;
                11'b000_0101_0011 : b_rgb<=1'b1;
                11'b000_0110_0011 : b_rgb<=1'b1;
                11'b000_0111_0011 : b_rgb<=1'b1;
                11'b000_1000_0011 : b_rgb<=1'b1;
                11'b000_1001_0011 : b_rgb<=1'b1;
                11'b000_1010_0011 : b_rgb<=1'b1;

                11'b000_0100_0100 : b_rgb<=1'b1;
                11'b000_1011_0100 : b_rgb<=1'b1;

                11'b000_0100_0101 : b_rgb<=1'b1;
                11'b000_1011_0101 : b_rgb<=1'b1;

                11'b000_0100_0110 : b_rgb<=1'b1;
                11'b000_1011_0110 : b_rgb<=1'b1;

                11'b000_0100_0111 : b_rgb<=1'b1;
                11'b000_0101_0111 : b_rgb<=1'b1;
                11'b000_0110_0111 : b_rgb<=1'b1;
                11'b000_0111_0111 : b_rgb<=1'b1;
                11'b000_1000_0111 : b_rgb<=1'b1;
                11'b000_1001_0111 : b_rgb<=1'b1;
                11'b000_1010_0111 : b_rgb<=1'b1;

                11'b000_0100_1000 : b_rgb<=1'b1;

                11'b000_0100_1001 : b_rgb<=1'b1;

                11'b000_0100_1010 : b_rgb<=1'b1;

                11'b000_0100_1011 : b_rgb<=1'b1;

                11'b000_0100_1100 : b_rgb<=1'b1;


                // A character

                11'b001_0100_0011 : b_rgb<=1'b1;
                11'b001_0101_0011 : b_rgb<=1'b1;
                11'b001_0110_0011 : b_rgb<=1'b1;
                11'b001_0111_0011 : b_rgb<=1'b1;
                11'b001_1000_0011 : b_rgb<=1'b1;
                11'b001_1001_0011 : b_rgb<=1'b1;
                11'b001_1010_0011 : b_rgb<=1'b1;
                11'b001_1011_0011 : b_rgb<=1'b1;

                11'b001_0100_0100 : b_rgb<=1'b1;
                11'b001_1011_0100 : b_rgb<=1'b1;

                11'b001_0100_0101 : b_rgb<=1'b1;
                11'b001_1011_0101 : b_rgb<=1'b1;

                11'b001_0100_0110 : b_rgb<=1'b1;
                11'b001_1011_0110 : b_rgb<=1'b1;

                11'b001_0100_0111 : b_rgb<=1'b1;
                11'b001_0101_0111 : b_rgb<=1'b1;
                11'b001_0110_0111 : b_rgb<=1'b1;
                11'b001_0111_0111 : b_rgb<=1'b1;
                11'b001_1000_0111 : b_rgb<=1'b1;
                11'b001_1001_0111 : b_rgb<=1'b1;
                11'b001_1010_0111 : b_rgb<=1'b1;
                11'b001_1011_0111 : b_rgb<=1'b1;

                11'b001_0100_1000 : b_rgb<=1'b1;
                11'b001_1011_1000 : b_rgb<=1'b1;

                11'b001_0100_1001 : b_rgb<=1'b1;
                11'b001_1011_1001 : b_rgb<=1'b1;

                11'b001_0100_1010 : b_rgb<=1'b1;
                11'b001_1011_1010 : b_rgb<=1'b1;

                11'b001_0100_1011 : b_rgb<=1'b1;
                11'b001_1011_1011 : b_rgb<=1'b1;

                11'b001_0100_1100 : b_rgb<=1'b1;
                11'b001_1011_1100 : b_rgb<=1'b1;

                // U character

                11'b010_0100_0011 : b_rgb<=1'b1;
                11'b010_1011_0011 : b_rgb<=1'b1;

                11'b010_0100_0100 : b_rgb<=1'b1;
                11'b010_1011_0100 : b_rgb<=1'b1;

                11'b010_0100_0101 : b_rgb<=1'b1;
                11'b010_1011_0101 : b_rgb<=1'b1;

                11'b010_0100_0110 : b_rgb<=1'b1;
                11'b010_1011_0110 : b_rgb<=1'b1;

                11'b010_0100_0111 : b_rgb<=1'b1;
                11'b010_1011_0111 : b_rgb<=1'b1;
                
                11'b010_0100_1000 : b_rgb<=1'b1;
                11'b010_1011_1000 : b_rgb<=1'b1;
                
                11'b010_0100_1001 : b_rgb<=1'b1;
                11'b010_1011_1001 : b_rgb<=1'b1;

                11'b010_0100_1010 : b_rgb<=1'b1;
                11'b010_1011_1010 : b_rgb<=1'b1;

                11'b010_0100_1011 : b_rgb<=1'b1;
                11'b010_1011_1011 : b_rgb<=1'b1;

                11'b010_0101_1100 : b_rgb<=1'b1;
                11'b010_0110_1100 : b_rgb<=1'b1;
                11'b010_0111_1100 : b_rgb<=1'b1;
                11'b010_1000_1100 : b_rgb<=1'b1;
                11'b010_1001_1100 : b_rgb<=1'b1;
                11'b010_1010_1100 : b_rgb<=1'b1;

                // S character

                11'b011_0100_0011 : b_rgb<=1'b1;
                11'b011_0101_0011 : b_rgb<=1'b1;
                11'b011_0110_0011 : b_rgb<=1'b1;
                11'b011_0111_0011 : b_rgb<=1'b1;
                11'b011_1000_0011 : b_rgb<=1'b1;
                11'b011_1001_0011 : b_rgb<=1'b1;
                11'b011_1010_0011 : b_rgb<=1'b1;
                11'b011_1011_0011 : b_rgb<=1'b1;

                11'b011_0100_0100 : b_rgb<=1'b1;

                11'b011_0100_0101 : b_rgb<=1'b1;

                11'b011_0100_0110 : b_rgb<=1'b1;

                11'b011_0100_0111 : b_rgb<=1'b1;
                11'b011_0101_0111 : b_rgb<=1'b1;
                11'b011_0110_0111 : b_rgb<=1'b1;
                11'b011_0111_0111 : b_rgb<=1'b1;
                11'b011_1000_0111 : b_rgb<=1'b1;
                11'b011_1001_0111 : b_rgb<=1'b1;
                11'b011_1010_0111 : b_rgb<=1'b1;
                11'b011_1011_0111 : b_rgb<=1'b1;

                11'b011_1011_1000 : b_rgb<=1'b1;

                11'b011_1011_1001 : b_rgb<=1'b1;

                11'b011_1011_1010 : b_rgb<=1'b1;

                11'b011_1011_1011 : b_rgb<=1'b1;

                11'b011_0100_1100 : b_rgb<=1'b1;
                11'b011_0101_1100 : b_rgb<=1'b1;
                11'b011_0110_1100 : b_rgb<=1'b1;
                11'b011_0111_1100 : b_rgb<=1'b1;
                11'b011_1000_1100 : b_rgb<=1'b1;
                11'b011_1001_1100 : b_rgb<=1'b1;
                11'b011_1010_1100 : b_rgb<=1'b1;
                11'b011_1011_1100 : b_rgb<=1'b1;

                // E character

                11'b100_0100_0011 : b_rgb<=1'b1;
                11'b100_0101_0011 : b_rgb<=1'b1;
                11'b100_0110_0011 : b_rgb<=1'b1;
                11'b100_0111_0011 : b_rgb<=1'b1;
                11'b100_1000_0011 : b_rgb<=1'b1;
                11'b100_1001_0011 : b_rgb<=1'b1;
                11'b100_1010_0011 : b_rgb<=1'b1;
                11'b100_1011_0011 : b_rgb<=1'b1;

                11'b100_0100_0100 : b_rgb<=1'b1;

                11'b100_0100_0101 : b_rgb<=1'b1;

                11'b100_0100_0110 : b_rgb<=1'b1;

                11'b100_0100_0111 : b_rgb<=1'b1;
                11'b100_0101_0111 : b_rgb<=1'b1;
                11'b100_0110_0111 : b_rgb<=1'b1;
                11'b100_0111_0111 : b_rgb<=1'b1;
                11'b100_1000_0111 : b_rgb<=1'b1;
                11'b100_1001_0111 : b_rgb<=1'b1;
                11'b100_1010_0111 : b_rgb<=1'b1;
                11'b100_1011_0111 : b_rgb<=1'b1;

                11'b100_0100_1000 : b_rgb<=1'b1;

                11'b100_0100_1001 : b_rgb<=1'b1;

                11'b100_0100_1010 : b_rgb<=1'b1;

                11'b100_0100_1011 : b_rgb<=1'b1;

                11'b100_0100_1100 : b_rgb<=1'b1;
                11'b100_0101_1100 : b_rgb<=1'b1;
                11'b100_0110_1100 : b_rgb<=1'b1;
                11'b100_0111_1100 : b_rgb<=1'b1;
                11'b100_1000_1100 : b_rgb<=1'b1;
                11'b100_1001_1100 : b_rgb<=1'b1;
                11'b100_1010_1100 : b_rgb<=1'b1;
                11'b100_1011_1100 : b_rgb<=1'b1;


                // D character

                11'b101_0100_0011 : b_rgb<=1'b1;
                11'b101_0101_0011 : b_rgb<=1'b1;
                11'b101_0110_0011 : b_rgb<=1'b1;
                11'b101_0111_0011 : b_rgb<=1'b1;
                11'b101_1000_0011 : b_rgb<=1'b1;
                11'b101_1001_0011 : b_rgb<=1'b1;

                11'b101_0100_0100 : b_rgb<=1'b1;
                11'b101_1010_0100 : b_rgb<=1'b1;

                11'b101_0100_0101 : b_rgb<=1'b1;
                11'b101_1011_0101 : b_rgb<=1'b1;

                11'b101_0100_0110 : b_rgb<=1'b1;
                11'b101_1011_0110 : b_rgb<=1'b1;

                11'b101_0100_0111 : b_rgb<=1'b1;
                11'b101_1011_0111 : b_rgb<=1'b1;

                11'b101_0100_1000 : b_rgb<=1'b1;
                11'b101_1011_1000 : b_rgb<=1'b1;

                11'b101_0100_1001 : b_rgb<=1'b1;
                11'b101_1011_1001 : b_rgb<=1'b1;

                11'b101_0100_1010 : b_rgb<=1'b1;
                11'b101_1011_1010 : b_rgb<=1'b1;

                11'b101_0100_1011 : b_rgb<=1'b1;
                11'b101_1010_1011 : b_rgb<=1'b1;

                11'b101_0100_1100 : b_rgb<=1'b1;
                11'b101_0101_1100 : b_rgb<=1'b1;
                11'b101_0110_1100 : b_rgb<=1'b1;
                11'b101_0111_1100 : b_rgb<=1'b1;
                11'b101_1000_1100 : b_rgb<=1'b1;
                11'b101_1001_1100 : b_rgb<=1'b1;



                default: b_rgb<=1'h0;
            endcase
            
        end


    assign pause_on = (pause) & (x>X_START & x<X_END & y>Y_START & y<Y_END) ? 1 :0;
    assign pause_rgb=b_rgb? 12'hfff :12'h000;

endmodule
